.CLK_50M_FPGA,
    .CLK_ENET_FPGA_P,
    .sw,
    .pb,
    .led,
    .mem_ck,
    .mem_ck_n,
    .mem_a,
    .mem_act_n,
    .mem_ba,
    .mem_bg,
    .mem_cke,
    .mem_cs_n,
    .mem_odt,
    .mem_reset_n,
    .mem_par,
    .mem_alert_n,
    .global_reset_reset_n,
    .pll_ref_clk,
    .oct_rzqin,
    .mem_dqs,
    .mem_dqs_n,
    .mem_dq,
    .mem_dbi_n,
    .pcie_perstn,
    .pcie_refclk,
    .pcie_rx,
    .pcie_tx,
    .user_led
